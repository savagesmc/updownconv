Upper VHF Bandpass Filter

V1 SRC 0 DC 0 AC 1 PULSE( 0 5 1u 1u 1u 1 1)
R1 SRC IN 50

C1 IN 0 30p
L1 IN 0 56n

C2 IN N2 13p
L2 N2 N3 130n

C3 N3 0 68p
L3 N3 0 24n

C4 N3 N4 10p
L4 N4 N5 160n

C5 N5 0 68p
L5 N5 0 24n

C6 N5 N6 10p
L6 N6 N7 160n

C7 N7 0 68p
L7 N7 0 24n

C8 N7 N8 13p
L8 N8 OUT 130n

C9 OUT 0 30p
L9 OUT 0 56n
R2 OUT 0 50

.control
   let mc_runs = 1000
   let run = 1
   set curplot = new
   set scratch = $curplot

   let tol = 0.01

   define unif(nom, var) (nom + nom*var * sunif(0))

   dowhile run <= mc_runs

      alter C1 = unif(30p, $tol)
      alter L1 = unif(56n, $tol)

      alter C2 = unif(13p, $tol)
      alter L2 = unif(130n, $tol)

      alter C3 = unif(68p, $tol)
      alter L3 = unif(24n, $tol)

      alter C4 = unif(10p, $tol)
      alter L4 = unif(160n, $tol)

      alter C5 = unif(68p, $tol)
      alter L5 = unif(24n, $tol)

      alter C6 = unif(10p, $tol)
      alter L6 = unif(160n, $tol)

      alter C7 = unif(68p, $tol)
      alter L7 = unif(24n, $tol)

      alter C8 = unif(13p, $tol)
      alter L8 = unif(130n, $tol)

      alter C9 = unif(30p, $tol)
      alter L9 = unif(56n, $tol)

      ac oct 100 10e6 500e6

      set run ="$&run"
      set dt = $curplot
      setplot $scratch

      let loss{$run}={$dt}.v(out)/{$dt}.v(in)
      setplot $dt
      let run = run + 1
   end
   set nolegend
   plot db({$scratch}.all) xlimit 50e6 300e6 ylimit -55 5 ylabel 'Upper VHF BPF - insertion loss'
.endc
.end
